`timescale 1ns/1ps

module simm (
  input 	   [17:0] addr,
  input 	   [1:0]ras,
  input 	   [3:0]cas,
  input		   we,
  output reg [15:0] data_out
);



endmodule
